module RAMfiller(
	input logic RAMsource,
	output logic RAMdata);
	
endmodule	